// module fp_add_sub(
//     input IEEE_extended_fp x1,
//     input IEEE_extended_fp x2,
//     input fp_op_t op,
//     input switched, //if the operands were switched during normalization
//     output IEEE_extended_fp ans
// )

// if(op == fp_add)


// endmodule