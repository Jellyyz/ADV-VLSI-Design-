// import fp_types::*; 

// module exponent_compare
// // take the exponents and compare them, and put out the result - may get more commplicated with more operations added
// (
//     input logic [7:0] exp1,
//     input logic [7:0] exp2,
//     input fp_op_t op
//     output logic [7:0] difference
// );


//     assign difference = exp1-exp2;

// endmodule