// //if systhesis tool is bad, we can optimize this, currently not using the module

// module twos_comp #(
//     parameter len = 22
// )
// (
//     input logic[len-1:0] in,
//     output logic[len-1:0] out
// );



// endmodule