module on_chip_sram

