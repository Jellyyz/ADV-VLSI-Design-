// import fp_types::*

// module flt_IEEE